module not1(a,c);
input a;
output c;
assign c=!a;
endmodule